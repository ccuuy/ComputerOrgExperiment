`timescale 1ns / 1ps

// 查找表乘法器实现
module mul4c(
	input clk,
	input[3:0] A,
	input[3:0] B,
	output reg[7:0]r
	);
	reg state = 0;
	reg [4:0]add;
	reg [4:0]sub;
	reg [7:0]a1;
	reg [7:0]b1;
    
	always @(posedge clk) begin
		if(state == 0)
		begin
			add = A + B;
			sub = A + (~B + 1);
			if (add[4] == 1)
				add = ~add + 1;
			if (sub[4] == 1)
				sub = ~sub + 1;
			state = state + 1;
		end
		else if(state == 1)
		begin
			case(add)
			5'b00000:a1 = 8'b00000000;
			5'b00001:a1 = 8'b00000000;
			5'b00010:a1 = 8'b00000001;
			5'b00011:a1 = 8'b00000010;
			5'b00100:a1 = 8'b00000100;
			5'b00101:a1 = 8'b00000110;
			5'b00110:a1 = 8'b00001001;
			5'b00111:a1 = 8'b00001100;
			5'b01000:a1 = 8'b00010000;
			5'b01001:a1 = 8'b00010100;
			5'b01010:a1 = 8'b00011001;
			5'b01011:a1 = 8'b00011110;
			5'b01100:a1 = 8'b00100100;
			5'b01101:a1 = 8'b00101010;
			5'b01110:a1 = 8'b00110001;
			5'b01111:a1 = 8'b00111000;
			endcase
			case(sub)
			5'b00000:b1 = 8'b00000000;
			5'b00001:b1 = 8'b00000000;
			5'b00010:b1 = 8'b00000001;
			5'b00011:b1 = 8'b00000010;
			5'b00100:b1 = 8'b00000100;
			5'b00101:b1 = 8'b00000110;
			5'b00110:b1 = 8'b00001001;
			5'b00111:b1 = 8'b00001100;
			5'b01000:b1 = 8'b00010000;
			5'b01001:b1 = 8'b00010100;
			5'b01010:b1 = 8'b00011001;
			5'b01011:b1 = 8'b00011110;
			5'b01100:b1 = 8'b00100100;
			5'b01101:b1 = 8'b00101010;
			5'b01110:b1 = 8'b00110001;
			5'b01111:b1 = 8'b00111000;
			endcase
			r = a1 + (~b1 + 1);
			state = state + 1;
		end

	end

endmodule
