module mult4(
 input [3:0] a, 
 input [3:0] b, 
 output [7:0] z , // 乘积输出 z
output ZF; // 标志位，不强制要求输出
 );
 
endmodule